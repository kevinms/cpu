module soc(

);
	
endmodule
